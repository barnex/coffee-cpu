module COFFEE(input CLK50);

wire address

module memory (
	address,
	clock,
	data,
	wren,
	q);
endmodule;
