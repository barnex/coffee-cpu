module COFFEE(input CLK50);

module memory (
	address,
	clock,
	data,
	wren,
	q);
endmodule;
